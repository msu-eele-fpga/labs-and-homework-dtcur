--Required packages
--Must be compiled with 2008 VHDL standard
library ieee;
use ieee.std_logic_1164.all;
-- Class packages
use work.print_pkg.all;
use work.assert_pkg.all;

